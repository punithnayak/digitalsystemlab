module program(a,f);
input a;
output f;
assign f= ~(~a);
endmodule	
